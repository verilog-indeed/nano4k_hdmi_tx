//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Device: GW1NSR-4C
//Created Time: Thu Sep 08 01:24:38 2022

module sp_framebuffer (dout, clk, oce, ce, reset, wre, ad, din);

output [5:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [14:0] ad;
input [5:0] din;

wire [30:0] sp_inst_0_dout_w;
wire [0:0] sp_inst_0_dout;
wire [30:0] sp_inst_1_dout_w;
wire [1:1] sp_inst_1_dout;
wire [29:0] sp_inst_2_dout_w;
wire [1:0] sp_inst_2_dout;
wire [30:0] sp_inst_3_dout_w;
wire [2:2] sp_inst_3_dout;
wire [30:0] sp_inst_4_dout_w;
wire [3:3] sp_inst_4_dout;
wire [29:0] sp_inst_5_dout_w;
wire [3:2] sp_inst_5_dout;
wire [30:0] sp_inst_6_dout_w;
wire [4:4] sp_inst_6_dout;
wire [30:0] sp_inst_7_dout_w;
wire [5:5] sp_inst_7_dout;
wire [29:0] sp_inst_8_dout_w;
wire [5:4] sp_inst_8_dout;
wire dff_q_0;
wire ce_w;
wire gw_gnd;

assign ce_w = ~wre & ce;
assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[30:0],sp_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 1;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_18 = 256'hEFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_19 = 256'h9F3DCF7F9F07FFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFF9F818F78FF1FFFFFFFF;
defparam sp_inst_0.INIT_RAM_1A = 256'h7FFFF800000FFFFFFFF9F3DE37F9F13FFFFFFFEFFFFFFFFFFFFC001FFFFFFFFF;
defparam sp_inst_0.INIT_RAM_1B = 256'hFFF1FFFCE33DEF711EF7FFFE0000003FFFFFFFDF3DFB7FCF1FFFE03C3E0FC5EF;
defparam sp_inst_0.INIT_RAM_1C = 256'h000003FFFFFFFFC1FD7C6F1FFFCF3BDEF7B9EF7FFF80000000FFFFFFFDFBDFD7;
defparam sp_inst_0.INIT_RAM_1D = 256'hFE300EF3BDEF7FFC000000001FFFFFFFF3DFC798F1FFFFE37EEFBBDEF7FFE000;
defparam sp_inst_0.INIT_RAM_1E = 256'hFFFFFFF7DFB77EF1FFFFE3FEEFBBDEF7FF00000000007FFFFFFF3DF977EF1FFF;
defparam sp_inst_0.INIT_RAM_1F = 256'h3BDE23FC00000000001FFFFFFFBDF377DF1FFFFE3FDE7BBDE73FC00000000001;
defparam sp_inst_0.INIT_RAM_20 = 256'hC1DF7C3C07FFFE303ECFBDE87F800000000000FFFFF9F1DCF71DF1FFFFE3FCE2;
defparam sp_inst_0.INIT_RAM_21 = 256'h0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFF9F;
defparam sp_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sp_inst_0.INIT_RAM_23 = 256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFF001FFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000F83E0;
defparam sp_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFE600000003FFFFFFFFFFFFFFFFFFF;
defparam sp_inst_0.INIT_RAM_26 = 256'hFFFC001F80700000001FFFFFFFF8000000000000000FFFFFC001FC0600000001;
defparam sp_inst_0.INIT_RAM_27 = 256'hF8000000000000000FFFFF8001F00300000000FFFFFFFF8000000000000000FF;
defparam sp_inst_0.INIT_RAM_28 = 256'h0003800000007FFFFFFF8000000000000000FFFFF8000000300000000FFFFFFF;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000FFFFF00000001800000007FFFFFFF8000000000000000FFFFF0000;
defparam sp_inst_0.INIT_RAM_2A = 256'h000003FFFFFFF8000000000000000FFFFE00000003800000003FFFFFFF800000;
defparam sp_inst_0.INIT_RAM_2B = 256'hF7FFFFFE00000001800000003FFFFFFF8000000000000000FFFFE00000001800;
defparam sp_inst_0.INIT_RAM_2C = 256'hFFFFFFFF7F7F7F7F7F7F7FFFFFE00000001A00000003FFFFFFFFF7F7F7F7F7F7;
defparam sp_inst_0.INIT_RAM_2D = 256'hC000003FFFFC000001FFFFFFFFF7F7F7F7F7F7F7FFFFFE0000007FFE0000003F;
defparam sp_inst_0.INIT_RAM_2E = 256'hF7F7F7F7F7F7F7FFFFFC000007FFFFF850001FFFFFFFFF7F7F7F7F7F7F7FFFFF;
defparam sp_inst_0.INIT_RAM_2F = 256'hFFFFFFFC001FFFFFFFFF7F7F7F7F7F7F7FFFFFC001F9FFFFFFCF8001FFFFFFFF;
defparam sp_inst_0.INIT_RAM_30 = 256'h00000000FFFFC003FFFFFFFFFFE001FFFFFFFFF7F7F7F7F7F7F7FFFFFC003FFF;
defparam sp_inst_0.INIT_RAM_31 = 256'hE001FFFFFFFC000000000000001FFFFC003FFFFFFFFFFF001FFFFFFF80000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h1FFFFC003FFC1FFC1FFF001FFFFFFFC000000000000001FFFFC007FFF7FFF7FF;
defparam sp_inst_0.INIT_RAM_33 = 256'hFFFFC000000000000001FFFFC003FFC1FFC0FFE001FFFFFFFC00000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h01FF80FF80FF8001FFFFFFFC000000000000001FFFFC003FF80FF80FFC001FFF;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000001FFFFC000FF80FFC0FF8001FFFFFFFC000000000000001FFFFC0;
defparam sp_inst_0.INIT_RAM_36 = 256'hFF7FF0003FFFFFFF8000000000000000FFFFC000FFC1FFC1FF8001FFFFFFFC00;
defparam sp_inst_0.INIT_RAM_37 = 256'h7F7F7EFFFFE000FFFFFFFFFF8003FFFFFFFBF7F7F7F7F7F7F7EFFFFE000FFF3F;
defparam sp_inst_0.INIT_RAM_38 = 256'h03FFFFFFFBF7F7F7F7F7F7F7EFFFFE000FFFFFFFFFF0003FFFFFFFBF7F7F7F7F;
defparam sp_inst_0.INIT_RAM_39 = 256'hFFFE0003FFFFFFFFE0003FFFFFFFBF7F7F7F7F7F7F7EFFFFE0007FFFFFFFFF00;
defparam sp_inst_0.INIT_RAM_3A = 256'hFFBF7F7F7F7F7F7F7EFFFFF0003FF7FFE7FE0007FFFFFFFBF7F7F7F7F7F7F7EF;
defparam sp_inst_0.INIT_RAM_3B = 256'h1FFC1C1FF8000FFFFFFFFBF7F7F7F7F7F7F7EFFFFF0001FF0FFC7FC0007FFFFF;
defparam sp_inst_0.INIT_RAM_3C = 256'h00000000000FFFFF8000FFE003FF0000FFFFFFFF8000000000000000FFFFF800;
defparam sp_inst_0.INIT_RAM_3D = 256'hFC0001FFFFFFFF8000000000000000FFFFFC0003FFFFFFE0001FFFFFFFF80000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000FFFFFE00003FFFFF00003FFFFFFFF8000000000000000FFFFFC0000FFFFF;
defparam sp_inst_0.INIT_RAM_3F = 256'hFFFFFFF8000000000000000FFFFFF000007FFF000007FFFFFFFF800000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[30:0],sp_inst_1_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 1;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_18 = 256'hCFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_19 = 256'h9F9CE73F3FA7FFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF9FC0CF387F9FFFFFFFF;
defparam sp_inst_1.INIT_RAM_1A = 256'h3FFFFC00001FFFFFFFF9FBCF73FDFBBFFFFFFFCFFFFFFFFFFFF8000FFFFFFFFF;
defparam sp_inst_1.INIT_RAM_1B = 256'hFCFBFFFCC799CE7B8CF3FFFE0000003FFFFFFF9FBCF33FDFBFFFE37C3C0F84CF;
defparam sp_inst_1.INIT_RAM_1C = 256'h000003FFFFFF9FC0FC380FBFFFDE73CCF33CCF3FFF80000000FFFFFFF9F9CF93;
defparam sp_inst_1.INIT_RAM_1D = 256'hFF700CFB3CCF3FF8000000000FFFFFF9F9CFC33CFBFFFFF73CCF33CCF3FFE000;
defparam sp_inst_1.INIT_RAM_1E = 256'hFFFFF9F3CF333CFBFFFFF7FCCF33CCF3FF00000000007FFFFF9F3CF933CFBFFF;
defparam sp_inst_1.INIT_RAM_1F = 256'h73CC77F800000000000FFFFFFF3CE733CFBFFFFF7FCCF33CCF7FE00000000003;
defparam sp_inst_1.INIT_RAM_20 = 256'hC08F3C3C03FFFF783C873CC8FF0000000000007FFFF9FBCE73B9FBFFFFF7F9C7;
defparam sp_inst_1.INIT_RAM_21 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000003FFFF9F;
defparam sp_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sp_inst_1.INIT_RAM_23 = 256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_24 = 256'hFFFFFFFFFFE001FFFE00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000F07E0;
defparam sp_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFC600000003FFFFFFFFFFFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_26 = 256'hFFFC001F80300000001FFFFFFFF8000000000000000FFFFFC001FC0700000001;
defparam sp_inst_1.INIT_RAM_27 = 256'hF8000000000000000FFFFF8000F80300000000FFFFFFFF8000000000000000FF;
defparam sp_inst_1.INIT_RAM_28 = 256'h0003000000007FFFFFFF8000000000000000FFFFF8000600300000000FFFFFFF;
defparam sp_inst_1.INIT_RAM_29 = 256'h0000000000FFFFF00000003800000007FFFFFFF8000000000000000FFFFF0000;
defparam sp_inst_1.INIT_RAM_2A = 256'h000003FFFFFFF8000000000000000FFFFF00000001800000007FFFFFFF800000;
defparam sp_inst_1.INIT_RAM_2B = 256'h000FFFFE00000001800000003FFFFFFF8000000000000000FFFFE00000001800;
defparam sp_inst_1.INIT_RAM_2C = 256'hFFFFFF8000000000000000FFFFE00000001C00000003FFFFFFF8000000000000;
defparam sp_inst_1.INIT_RAM_2D = 256'hC000001FFFFE000001FFFFFFF8000000000000000FFFFC0000003FFF0000001F;
defparam sp_inst_1.INIT_RAM_2E = 256'h000000000000000FFFFC00000FFFFFF820001FFFFFFF8000000000000000FFFF;
defparam sp_inst_1.INIT_RAM_2F = 256'hFFFFFFFE001FFFFFFF8000000000000000FFFFC000F9FFFFFFFFC001FFFFFFF8;
defparam sp_inst_1.INIT_RAM_30 = 256'h00000000FFFFC003FFFFFFFFFFE001FFFFFFF8000000000000000FFFFC001FFF;
defparam sp_inst_1.INIT_RAM_31 = 256'hF001FFFFFFFBF7F7F7F7F7F7F7EFFFFC007FFFFFFFFFFE001FFFFFFF80000000;
defparam sp_inst_1.INIT_RAM_32 = 256'hEFFFFC007FFC1FFC1FFE001FFFFFFFBF7F7F7F7F7F7F7EFFFFC007FFFFFFFFFF;
defparam sp_inst_1.INIT_RAM_33 = 256'hFFFFBF7F7F7F7F7F7F7EFFFFC003FF80FF80FFE001FFFFFFFBF7F7F7F7F7F7F7;
defparam sp_inst_1.INIT_RAM_34 = 256'h01FF80FF80FFC001FFFFFFFBF7F7F7F7F7F7F7EFFFFC003FF80FF80FFE001FFF;
defparam sp_inst_1.INIT_RAM_35 = 256'hF7F7F7F7F7F7EFFFFC000FF80FF80FF8001FFFFFFFBF7F7F7F7F7F7F7EFFFFC0;
defparam sp_inst_1.INIT_RAM_36 = 256'hFFFFF8001FFFFFFF8000000000000000FFFFC000FFC1FFC1FF8001FFFFFFFBF7;
defparam sp_inst_1.INIT_RAM_37 = 256'h7F7F7FFFFFE000FFFFFFFFFF0003FFFFFFFFF7F7F7F7F7F7F7FFFFFC000FFE7F;
defparam sp_inst_1.INIT_RAM_38 = 256'h03FFFFFFFFF7F7F7F7F7F7F7FFFFFE0007FFFFFFFFF0003FFFFFFFFF7F7F7F7F;
defparam sp_inst_1.INIT_RAM_39 = 256'hFFFF0007FFFFFFFFE0007FFFFFFFFF7F7F7F7F7F7F7FFFFFE0007FFFFFFFFF00;
defparam sp_inst_1.INIT_RAM_3A = 256'hFFFF7F7F7F7F7F7F7FFFFFF0003FF3FFE7FE0007FFFFFFFFF7F7F7F7F7F7F7FF;
defparam sp_inst_1.INIT_RAM_3B = 256'h0FF8000FF8000FFFFFFFFFF7F7F7F7F7F7F7FFFFFF0001FF1FF87FC0007FFFFF;
defparam sp_inst_1.INIT_RAM_3C = 256'h00000000000FFFFF80007FF007FF0000FFFFFFFF8000000000000000FFFFF800;
defparam sp_inst_1.INIT_RAM_3D = 256'hF80001FFFFFFFF8000000000000000FFFFFC0003FFFFFFE0001FFFFFFFF80000;
defparam sp_inst_1.INIT_RAM_3E = 256'h0000FFFFFE00007FFFFE00003FFFFFFFF8000000000000000FFFFFC0001FFFFF;
defparam sp_inst_1.INIT_RAM_3F = 256'hFFFFFFF8000000000000000FFFFFE00000FFFF800003FFFFFFFF800000000000;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[29:0],sp_inst_2_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b00;
defparam sp_inst_2.BIT_WIDTH = 2;
defparam sp_inst_2.BLK_SEL = 3'b010;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'h00000000000000000000FFFFFFFFFFFF0000000000006FFE4000000000003FFF;
defparam sp_inst_2.INIT_RAM_01 = 256'hFFFFFFC000000000000000000000000000FFFFFFFFFFFFFFFFFFC00000000000;
defparam sp_inst_2.INIT_RAM_02 = 256'h00000002FFFFFFFFFFFFFFFFFFC0000000000000000000000000000000FFFFFF;
defparam sp_inst_2.INIT_RAM_03 = 256'hC0000000000000000000000000000000FFFFFFFFFFFFE0000000000000000000;
defparam sp_inst_2.INIT_RAM_04 = 256'h551555FFFFFFFFFFFFF400000000000000000000000007FFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_05 = 256'h0000000000000000001FFFFFFFFFFFFFFFFFFFD5551555155515551555155515;
defparam sp_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFD5551555155515551555155515551555FFFFFFFFFFFFFD000000;
defparam sp_inst_2.INIT_RAM_07 = 256'h551555155515551555FFFFFFFFFFFFFF4000000000000000000000007FFFFFFF;
defparam sp_inst_2.INIT_RAM_08 = 256'hFFFFFFD00000000000000000000001FFFFFFFFFFFFFFFFFFFFD5551555155515;
defparam sp_inst_2.INIT_RAM_09 = 256'h000BFFFFFFFFFFFFFFFFFFFFD5551555155515551555155515551555FFFFFFFF;
defparam sp_inst_2.INIT_RAM_0A = 256'h551555155515551555155515551555FFFFFFFFFFFFFFF8000000000000000000;
defparam sp_inst_2.INIT_RAM_0B = 256'h1555FFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFFFD5;
defparam sp_inst_2.INIT_RAM_0C = 256'h00000000000001FFFFFFFFFFFFFFFFFFFFFFD555155515551555155515551555;
defparam sp_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFD5551555155515551555155515551555FFFFFFFFFFFFFFFFD00000;
defparam sp_inst_2.INIT_RAM_0E = 256'h0000000000000000FFFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_0F = 256'hFFFFFFFFC000000000000000FFFFFFFFFFFFFFFFFFFFFFFFC000000000000000;
defparam sp_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFDAAA2AAA2AAA2AAA2AAA2AAA2AAA2AA9FFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_11 = 256'h2AAA2AAA2AAA2AAA2AAA2AAA2AA9FFFFFFFFFFFFFFFFFFFC0000000000000FFF;
defparam sp_inst_2.INIT_RAM_12 = 256'hA9FFFFFFFFFFFFFFFFFFFFE00000000002FFFFFFFFFFFFFFFFFFFFFFFFFFDAAA;
defparam sp_inst_2.INIT_RAM_13 = 256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAA2AAA2AAA2AAA2AAA2AAA2AAA2A;
defparam sp_inst_2.INIT_RAM_14 = 256'hFFFFFFFFDAAA2AAA2AAA2AAA2AAA2AAA2AAA2AA9FFFFFFFFFFFFFFFFFFFFFFD0;
defparam sp_inst_2.INIT_RAM_15 = 256'hAA2AAA2AAA2AA9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAA2AAA2AAA2AAA2A;
defparam sp_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFDAAA2AAA2AAA2AAA2AAA2AAA2AAA2AA9FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_18 = 256'hAA2AAA2AAA2AAA2AAA2AAA2AA9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAA2A;
defparam sp_inst_2.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_1B = 256'hFFFFFFEFFF3FFF3FFF3FFF3FFF3FFF3FFF3FFEFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1C = 256'h3FFF3FFF3FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF3FFF3FFF3FFF;
defparam sp_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFEFFF3FFF3FFF3FFF3FFF3FFF3FFF3FFEFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1F = 256'h3FFF3FFF3FFF3FFF3FFF3FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF;
defparam sp_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF3FFF3FFF3FFF3FFF3FFF3FFEFF;
defparam sp_inst_2.INIT_RAM_22 = 256'hFFFFEFFF3FFF3FFF3FFF3FFF3FFF3FFF3FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_23 = 256'hAA2AAA2AA9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAA2AAA2AAA2AAA2AAA2A;
defparam sp_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_28 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[30:0],sp_inst_3_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b00;
defparam sp_inst_3.BIT_WIDTH = 1;
defparam sp_inst_3.BLK_SEL = 3'b000;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_05 = 256'h3FFFFFFFFFFF3FFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFCFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_07 = 256'hFF01FCFFFFFF3FFFFFFFFC3FC1FF00E01FFFFF3FFFFFFFF83FDFFFFFF7FFFFFF;
defparam sp_inst_3.INIT_RAM_08 = 256'h7CF8FFDFFFFFFFFFFFFFFFCFEFFFFFFBFFFFFFFFE3F80FE00E01FFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_09 = 256'hF803FCFFFFFFFF99FFF1DF8FFDFC73F07BFEF03FFE3CFFC33F3FFFFFFFFC3FFE;
defparam sp_inst_3.INIT_RAM_0A = 256'hF3C3F1FBFEC7C7FE3F7FDE3FDFFFFFFFFDDFFFB9F8FFDF813F07BFEF01FFF7F3;
defparam sp_inst_3.INIT_RAM_0B = 256'hFFFFFFF1CF870DF8F01E3E3F1F3DE6FEF0E1F3FCF3FCFFFFFFFF89FFF1DF8FFD;
defparam sp_inst_3.INIT_RAM_0C = 256'h98CC7C73E1F3FFFBFCFFFFFFFFBEF878878F01E3E3F1FBDEEFC70F1FBF8FBFEF;
defparam sp_inst_3.INIT_RAM_0D = 256'h3E79F0F80FFDE3E3F1FD25C7C73E1FCFFFBFF3FFFFFFF1CF9F0C00FFDE3E3F1F;
defparam sp_inst_3.INIT_RAM_0E = 256'h3C7FCFFFBFF3FFFFFFF0079F9FF8FFDE3E3F1FCB9EFC73F3FDFFFBFF7FFFFFFE;
defparam sp_inst_3.INIT_RAM_0F = 256'hF8FFDE3E3F1FD25E7C73C7FEFFFBFFBFFFFFFE0079E3FF8FFDE3E3F1FC71EFEF;
defparam sp_inst_3.INIT_RAM_10 = 256'hFBFFCFFFFFFEFFB807FF8FFDE3E3803870E01F00FFCFFFBFF3FFFFFFC7F39E3F;
defparam sp_inst_3.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFF7FFFFFDFFFFFFCFFBC1FFF8FFDE3E3803CF9FC1F83FFF3F;
defparam sp_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFCFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFEFF;
defparam sp_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_18 = 256'hEFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_19 = 256'h9F3DCF7F9F07FFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFF9F818F78FF1FFFFFFFF;
defparam sp_inst_3.INIT_RAM_1A = 256'h7FFFFBFFFFEFFFFFFFF9F3DE37F9F13FFFFFFFEFFFFFFFFFFFFBFFEFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_1B = 256'hFFF1FFFCE33DEF711EF7FFFFFFFFFFFFFFFFFFDF3DFB7FCF1FFFE03C3E0FC5EF;
defparam sp_inst_3.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFC1FD7C6F1FFFCF3BDEF7B9EF7FFFFFFFFFFFFFFFFFFDFBDFD7;
defparam sp_inst_3.INIT_RAM_1D = 256'hFE300EF3BDEF7FFBFFFFFFFFEFFFFFFFF3DFC798F1FFFFE37EEFBBDEF7FFFFFF;
defparam sp_inst_3.INIT_RAM_1E = 256'hFFFFFFF7DFB77EF1FFFFE3FEEFBBDEF7FFFFFFFFFFFFFFFFFFFF3DF977EF1FFF;
defparam sp_inst_3.INIT_RAM_1F = 256'h3BDE23FBFFFFFFFFFFEFFFFFFFBDF377DF1FFFFE3FDE7BBDE73FFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_20 = 256'hC1DF7C3C07FFFE303ECFBDE87FFFFFFFFFFFFFFFFFF9F1DCF71DF1FFFFE3FCE2;
defparam sp_inst_3.INIT_RAM_21 = 256'hFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9F;
defparam sp_inst_3.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD;
defparam sp_inst_3.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_24 = 256'hFFFFFFFFFFEFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF;
defparam sp_inst_3.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007F007F007F00FFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_27 = 256'hFC000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000FF;
defparam sp_inst_3.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFC000000000000000FFFFFFFFF9FFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_29 = 256'h0000000000FFFFFFFFFFFFDFFFFFFFFFFFFFFFFC000000000000000FFFFFFFFF;
defparam sp_inst_3.INIT_RAM_2A = 256'hFFFFFFFFFFFFFC000000000000000FFFFEFFFFFFFFFFFFFFFFBFFFFFFFC00000;
defparam sp_inst_3.INIT_RAM_2B = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_2C = 256'hFFFFFFC000000000000000FFFFFFFFFFFFFBFFFFFFFFFFFFFFFC000000000000;
defparam sp_inst_3.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000FFFFDFFFFFFFFFFFFFFFFDF;
defparam sp_inst_3.INIT_RAM_2E = 256'h000000000000000FFFFFFFFFF7FFFFFFCFFFFFFFFFFFC000000000000000FFFF;
defparam sp_inst_3.INIT_RAM_2F = 256'hFFFFFFFDFFFFFFFFFFC000000000000000FFFFFFFEFFFFFFFFCFBFFFFFFFFFFC;
defparam sp_inst_3.INIT_RAM_30 = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000FFFFFFFDFFF;
defparam sp_inst_3.INIT_RAM_31 = 256'hEFFFFFFFFFFC000000000000000FFFFFFFBFFFFFFFFFFEFFFFFFFFFF80000000;
defparam sp_inst_3.INIT_RAM_32 = 256'h0FFFFFFFBFFFFFFFFFFEFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFF7FF;
defparam sp_inst_3.INIT_RAM_33 = 256'hFFFFC000000000000000FFFFFFFFFFBFFFBFFFFFFFFFFFFFFC00000000000000;
defparam sp_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFBFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_35 = 256'h0000000000000FFFFFFFFFFFFFFBFFFFFFFFFFFFFFC000000000000000FFFFFF;
defparam sp_inst_3.INIT_RAM_36 = 256'hFF7FF7FFDFFFFFFF8000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sp_inst_3.INIT_RAM_37 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000FFFFDFFFFFEBF;
defparam sp_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFC000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000;
defparam sp_inst_3.INIT_RAM_39 = 256'hFFFEFFFBFFFFFFFFFFFFBFFFFFFFC000000000000000FFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_3A = 256'hFFC000000000000000FFFFFFFFFFFBFFFFFFFFFFFFFFFFFC000000000000000F;
defparam sp_inst_3.INIT_RAM_3B = 256'hFFFBFFEFFFFFFFFFFFFFFC000000000000000FFFFFFFFFFFEFFBFFFFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_3C = 256'hF7F7F7F7F7FFFFFFFFFFFFEFFBFFFFFFFFFFFFFF8000000000000000FFFFFFFF;
defparam sp_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFBF7F7F7F7F7F7F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F7;
defparam sp_inst_3.INIT_RAM_3E = 256'h7F7FFFFFFFFFFFBFFFFFFFFFFFFFFFFFFBF7F7F7F7F7F7F7FFFFFFFFFFEFFFFF;
defparam sp_inst_3.INIT_RAM_3F = 256'hFFFFFFFBF7F7F7F7F7F7F7FFFFFFEFFFFFFFFF7FFFFBFFFFFFFFBF7F7F7F7F7F;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[30:0],sp_inst_4_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b00;
defparam sp_inst_4.BIT_WIDTH = 1;
defparam sp_inst_4.BLK_SEL = 3'b000;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_05 = 256'h1FFFFFFFFFFF9FFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFF9FFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_07 = 256'hFE00FCFFFFFF3FFFFFFFFE3F81FF01E00FFFFF1FFFFFFFF03F8FFFFFE3FFFFFF;
defparam sp_inst_4.INIT_RAM_08 = 256'h3879FF8FFFFFFFFFFFFFE787C7FFFFF1FFFFFFFFC1F007C01E00FFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_09 = 256'hFC09F9FFFFFFFFC9FFE38F9FF8F827F031FC783FFC7E7FE19F9FFFFFFFFC9F3C;
defparam sp_inst_4.INIT_RAM_0A = 256'hF187F3F1FC638FFF3E3F8C1F8FFFFFFFF88FFF18F9FF8F007F031FC600FFE3E7;
defparam sp_inst_4.INIT_RAM_0B = 256'hFFFFFFF9CF0398F9E00F3C7F3F98CC7C6073F3F9E1FCFFFFFFFF9CFFF98F9FF8;
defparam sp_inst_4.INIT_RAM_0C = 256'h98CCFE67F3F9FFF1FE7FFFFFFF1C7039C79E00F3E7F3F98CC7E6073F1F9F1FC7;
defparam sp_inst_4.INIT_RAM_0D = 256'h3E73F9F01FF8F3E7F3F98CCFE67F3F9FFF1FE7FFFFFFF3E73F9E01FF8F3E7F3F;
defparam sp_inst_4.INIT_RAM_0E = 256'h7E3FCFFF1FF3FFFFFFE0033F1FF9FF8F3E7F3F924C7E67E3F8FFF1FE3FFFFFFF;
defparam sp_inst_4.INIT_RAM_0F = 256'hF9FF8F3E7F3F870E38E787FC7FF1FF1FFFFFFE0033F1FF9FF8F3E7F3F924C7C6;
defparam sp_inst_4.INIT_RAM_10 = 256'hF1FF9FFFFFFC7F1007FF9FF8F3E7003C71F00E00FFE7FF1FF9FFFFFFE7F33C3F;
defparam sp_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFE3FFFFF8FFFFFFC7F180FFF9FF8F3E7003C71F83F01FFE7F;
defparam sp_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFCFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFC7F;
defparam sp_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_18 = 256'hCFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_19 = 256'h9F9CE73F3FA7FFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF9FC0CF387F9FFFFFFFF;
defparam sp_inst_4.INIT_RAM_1A = 256'h3FFFFC00001FFFFFFFF9FBCF73FDFBBFFFFFFFCFFFFFFFFFFFFC001FFFFFFFFF;
defparam sp_inst_4.INIT_RAM_1B = 256'hFCFBFFFCC799CE7B8CF3FFFE0000003FFFFFFF9FBCF33FDFBFFFE37C3C0F84CF;
defparam sp_inst_4.INIT_RAM_1C = 256'h000003FFFFFF9FC0FC380FBFFFDE73CCF33CCF3FFF80000000FFFFFFF9F9CF93;
defparam sp_inst_4.INIT_RAM_1D = 256'hFF700CFB3CCF3FFC000000001FFFFFF9F9CFC33CFBFFFFF73CCF33CCF3FFE000;
defparam sp_inst_4.INIT_RAM_1E = 256'hFFFFF9F3CF333CFBFFFFF7FCCF33CCF3FF00000000007FFFFF9F3CF933CFBFFF;
defparam sp_inst_4.INIT_RAM_1F = 256'h73CC77FC00000000001FFFFFFF3CE733CFBFFFFF7FCCF33CCF7FE00000000003;
defparam sp_inst_4.INIT_RAM_20 = 256'hC08F3C3C03FFFF783C873CC8FF0000000000007FFFF9FBCE73B9FBFFFFF7F9C7;
defparam sp_inst_4.INIT_RAM_21 = 256'h0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000003FFFF9F;
defparam sp_inst_4.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sp_inst_4.INIT_RAM_23 = 256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFF001FFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000F07E0;
defparam sp_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFC600000003FFFFFFFFFFFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_26 = 256'hFFFC001F80300000001FFFFFFFF8000000000000000FFFFFC001FC0700000001;
defparam sp_inst_4.INIT_RAM_27 = 256'hFBF007F007F007F00FFFFF8000F80300000000FFFFFFFFBF007F007F007F00FF;
defparam sp_inst_4.INIT_RAM_28 = 256'h0003000000007FFFFFFFBF007F007F007F00FFFFF8000600300000000FFFFFFF;
defparam sp_inst_4.INIT_RAM_29 = 256'h007F007F00FFFFF00000003800000007FFFFFFFBF007F007F007F00FFFFF0000;
defparam sp_inst_4.INIT_RAM_2A = 256'h000003FFFFFFFBF007F007F007F00FFFFF00000001800000007FFFFFFFBF007F;
defparam sp_inst_4.INIT_RAM_2B = 256'hF00FFFFE00000001800000003FFFFFFF8000000000000000FFFFE00000001800;
defparam sp_inst_4.INIT_RAM_2C = 256'hFFFFFFBF007F007F007F00FFFFE00000001C00000003FFFFFFFBF007F007F007;
defparam sp_inst_4.INIT_RAM_2D = 256'hC000001FFFFE000001FFFFFFFBF007F007F007F00FFFFE0000003FFF0000003F;
defparam sp_inst_4.INIT_RAM_2E = 256'hF007F007F007F00FFFFC00000FFFFFF830001FFFFFFFBF007F007F007F00FFFF;
defparam sp_inst_4.INIT_RAM_2F = 256'hFFFFFFFE001FFFFFFFBF007F007F007F00FFFFC001F9FFFFFFFFC001FFFFFFFB;
defparam sp_inst_4.INIT_RAM_30 = 256'h00000000FFFFC003FFFFFFFFFFE001FFFFFFFBF007F007F007F00FFFFC003FFF;
defparam sp_inst_4.INIT_RAM_31 = 256'hF001FFFFFFFBF007F007F007F00FFFFC007FFFFFFFFFFF001FFFFFFF80000000;
defparam sp_inst_4.INIT_RAM_32 = 256'h0FFFFC007FFC1FFC1FFF001FFFFFFFBF007F007F007F00FFFFC007FFFFFFFFFF;
defparam sp_inst_4.INIT_RAM_33 = 256'hFFFFBF007F007F007F00FFFFC003FFC0FFC0FFE001FFFFFFFBF007F007F007F0;
defparam sp_inst_4.INIT_RAM_34 = 256'h01FF80FF80FFC001FFFFFFFBF007F007F007F00FFFFC003FF80FF80FFE001FFF;
defparam sp_inst_4.INIT_RAM_35 = 256'h07F007F007F00FFFFC000FF80FFC0FF8001FFFFFFFBF007F007F007F00FFFFC0;
defparam sp_inst_4.INIT_RAM_36 = 256'hFFFFF8003FFFFFFF8000000000000000FFFFC000FFC1FFC1FF8001FFFFFFFBF0;
defparam sp_inst_4.INIT_RAM_37 = 256'h007F00FFFFE000FFFFFFFFFF0003FFFFFFFBF007F007F007F00FFFFE000FFF7F;
defparam sp_inst_4.INIT_RAM_38 = 256'h03FFFFFFFBF007F007F007F00FFFFE0007FFFFFFFFF0003FFFFFFFBF007F007F;
defparam sp_inst_4.INIT_RAM_39 = 256'hFFFF0007FFFFFFFFE0007FFFFFFFBF007F007F007F00FFFFE0007FFFFFFFFF00;
defparam sp_inst_4.INIT_RAM_3A = 256'hFFBF007F007F007F00FFFFF0003FF7FFE7FE0007FFFFFFFBF007F007F007F00F;
defparam sp_inst_4.INIT_RAM_3B = 256'h0FFC001FF8000FFFFFFFFBF007F007F007F00FFFFF0001FF1FFC7FC0007FFFFF;
defparam sp_inst_4.INIT_RAM_3C = 256'hF007F007F00FFFFF80007FF007FF0000FFFFFFFF8000000000000000FFFFF800;
defparam sp_inst_4.INIT_RAM_3D = 256'hF80001FFFFFFFFFF007F007F007F00FFFFFC0003FFFFFFE0001FFFFFFFFFF007;
defparam sp_inst_4.INIT_RAM_3E = 256'h7F00FFFFFE00007FFFFE00003FFFFFFFFFF007F007F007F00FFFFFC0001FFFFF;
defparam sp_inst_4.INIT_RAM_3F = 256'hFFFFFFFFF007F007F007F00FFFFFF00000FFFF800007FFFFFFFFFF007F007F00;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[29:0],sp_inst_5_dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b00;
defparam sp_inst_5.BIT_WIDTH = 2;
defparam sp_inst_5.BLK_SEL = 3'b010;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'h15553FFF15553FFF1555FFFFFFFFFFFF555555555555AFFE5555555555557FFF;
defparam sp_inst_5.INIT_RAM_01 = 256'hFFFFFFD555555555555555555555555555FFFFFFFFFFFFFFFFFFEFFF15553FFF;
defparam sp_inst_5.INIT_RAM_02 = 256'h55555557FFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFF;
defparam sp_inst_5.INIT_RAM_03 = 256'hC0000000000000000000000000000000FFFFFFFFFFFFF5555555555555555555;
defparam sp_inst_5.INIT_RAM_04 = 256'hFF1555FFFFFFFFFFFFF95555555555555555555555555BFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_05 = 256'h5555555555555555555FFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553F;
defparam sp_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFD555555;
defparam sp_inst_5.INIT_RAM_07 = 256'h553FFF15553FFF1555FFFFFFFFFFFFFF5555555555555555555555557FFFFFFF;
defparam sp_inst_5.INIT_RAM_08 = 256'hFFFFFFE55555555555555555555556FFFFFFFFFFFFFFFFFFFFEFFF15553FFF15;
defparam sp_inst_5.INIT_RAM_09 = 256'h555FFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFF;
defparam sp_inst_5.INIT_RAM_0A = 256'hFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFD555555555555555555;
defparam sp_inst_5.INIT_RAM_0B = 256'h1555FFFFFFFFFFFFFFFF555555555555555555557FFFFFFFFFFFFFFFFFFFFFEF;
defparam sp_inst_5.INIT_RAM_0C = 256'h55555555555556FFFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF;
defparam sp_inst_5.INIT_RAM_0D = 256'hFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFFE55555;
defparam sp_inst_5.INIT_RAM_0E = 256'h0000000000000000FFFFFFFFFFFFFFFFFD55555555555555555FFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_0F = 256'hFFFFFFFFD555555555555555FFFFFFFFFFFFFFFFFFFFFFFFC000000000000000;
defparam sp_inst_5.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_11 = 256'h15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFFFFFD5555555555555FFF;
defparam sp_inst_5.INIT_RAM_12 = 256'h55FFFFFFFFFFFFFFFFFFFFE55555555556FFFFFFFFFFFFFFFFFFFFFFFFFFEFFF;
defparam sp_inst_5.INIT_RAM_13 = 256'h555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF15;
defparam sp_inst_5.INIT_RAM_14 = 256'hFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFFFFFFFFE5;
defparam sp_inst_5.INIT_RAM_15 = 256'hFF15553FFF1555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553F;
defparam sp_inst_5.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_18 = 256'h553FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF15;
defparam sp_inst_5.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000;
defparam sp_inst_5.INIT_RAM_1B = 256'hFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_1C = 256'h15553FFF1555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF;
defparam sp_inst_5.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_1F = 256'h3FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF1555;
defparam sp_inst_5.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF15553FFF15553FFF15553FFF1555FF;
defparam sp_inst_5.INIT_RAM_22 = 256'hFFFFEFFF15553FFF15553FFF15553FFF1555FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_23 = 256'h552AAA1554FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAA15552AAA15552AAA15;
defparam sp_inst_5.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_5.INIT_RAM_28 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SP sp_inst_6 (
    .DO({sp_inst_6_dout_w[30:0],sp_inst_6_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]})
);

defparam sp_inst_6.READ_MODE = 1'b0;
defparam sp_inst_6.WRITE_MODE = 2'b00;
defparam sp_inst_6.BIT_WIDTH = 1;
defparam sp_inst_6.BLK_SEL = 3'b000;
defparam sp_inst_6.RESET_MODE = "SYNC";
defparam sp_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_18 = 256'hEFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_19 = 256'h9F3DCF7F9F07FFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFF9F818F78FF1FFFFFFFF;
defparam sp_inst_6.INIT_RAM_1A = 256'h7FFFFFFFFFFFFFFFFFF9F3DE37F9F13FFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_1B = 256'hFFF1FFFCE33DEF711EF7FFFFFFFFFFFFFFFFFFDF3DFB7FCF1FFFE03C3E0FC5EF;
defparam sp_inst_6.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFC1FD7C6F1FFFCF3BDEF7B9EF7FFFFFFFFFFFFFFFFFFDFBDFD7;
defparam sp_inst_6.INIT_RAM_1D = 256'hFE300EF3BDEF7FFFFFFFFFFFFFFFFFFFF3DFC798F1FFFFE37EEFBBDEF7FFFFFF;
defparam sp_inst_6.INIT_RAM_1E = 256'hFFFFFFF7DFB77EF1FFFFE3FEEFBBDEF7FFFFFFFFFFFFFFFFFFFF3DF977EF1FFF;
defparam sp_inst_6.INIT_RAM_1F = 256'h3BDE23FFFFFFFFFFFFFFFFFFFFBDF377DF1FFFFE3FDE7BBDE73FFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_20 = 256'hC1DF7C3C07FFFE303ECFBDE87FFFFFFFFFFFFFFFFFF9F1DCF71DF1FFFFE3FCE2;
defparam sp_inst_6.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9F;
defparam sp_inst_6.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007F7F7F7F0000FFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_27 = 256'hFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FF;
defparam sp_inst_6.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_29 = 256'h007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFF;
defparam sp_inst_6.INIT_RAM_2A = 256'hFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00;
defparam sp_inst_6.INIT_RAM_2B = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_2C = 256'hFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0;
defparam sp_inst_6.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_2E = 256'hF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFF;
defparam sp_inst_6.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFB;
defparam sp_inst_6.INIT_RAM_30 = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_31 = 256'hFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000;
defparam sp_inst_6.INIT_RAM_32 = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_33 = 256'hFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F000;
defparam sp_inst_6.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_35 = 256'hF00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFF;
defparam sp_inst_6.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7;
defparam sp_inst_6.INIT_RAM_37 = 256'h7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_38 = 256'hFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F;
defparam sp_inst_6.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_3A = 256'hFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000F;
defparam sp_inst_6.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_3C = 256'h0007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000FFFFFFFF;
defparam sp_inst_6.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F0;
defparam sp_inst_6.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFF;
defparam sp_inst_6.INIT_RAM_3F = 256'hFFFFFFFBF7F00007F7F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F00007F7F;

SP sp_inst_7 (
    .DO({sp_inst_7_dout_w[30:0],sp_inst_7_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]})
);

defparam sp_inst_7.READ_MODE = 1'b0;
defparam sp_inst_7.WRITE_MODE = 2'b00;
defparam sp_inst_7.BIT_WIDTH = 1;
defparam sp_inst_7.BLK_SEL = 3'b000;
defparam sp_inst_7.RESET_MODE = "SYNC";
defparam sp_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_18 = 256'hCFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_19 = 256'h9F9CE73F3FA7FFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF9FC0CF387F9FFFFFFFF;
defparam sp_inst_7.INIT_RAM_1A = 256'h3FFFFFFFFFFFFFFFFFF9FBCF73FDFBBFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_1B = 256'hFCFBFFFCC799CE7B8CF3FFFFFFFFFFFFFFFFFF9FBCF33FDFBFFFE37C3C0F84CF;
defparam sp_inst_7.INIT_RAM_1C = 256'hFFFFFFFFFFFF9FC0FC380FBFFFDE73CCF33CCF3FFFFFFFFFFFFFFFFFF9F9CF93;
defparam sp_inst_7.INIT_RAM_1D = 256'hFF700CFB3CCF3FFFFFFFFFFFFFFFFFF9F9CFC33CFBFFFFF73CCF33CCF3FFFFFF;
defparam sp_inst_7.INIT_RAM_1E = 256'hFFFFF9F3CF333CFBFFFFF7FCCF33CCF3FFFFFFFFFFFFFFFFFF9F3CF933CFBFFF;
defparam sp_inst_7.INIT_RAM_1F = 256'h73CC77FFFFFFFFFFFFFFFFFFFF3CE733CFBFFFFF7FCCF33CCF7FFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_20 = 256'hC08F3C3C03FFFF783C873CC8FFFFFFFFFFFFFFFFFFF9FBCE73B9FBFFFFF7F9C7;
defparam sp_inst_7.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9F;
defparam sp_inst_7.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFBF7F000000000000FFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_27 = 256'hFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FF;
defparam sp_inst_7.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_29 = 256'h7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFF;
defparam sp_inst_7.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F;
defparam sp_inst_7.INIT_RAM_2B = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_2C = 256'hFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000;
defparam sp_inst_7.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_2E = 256'hF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFF;
defparam sp_inst_7.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_30 = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_31 = 256'hFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000;
defparam sp_inst_7.INIT_RAM_32 = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_33 = 256'hFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F0000000;
defparam sp_inst_7.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_35 = 256'hF7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFF;
defparam sp_inst_7.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam sp_inst_7.INIT_RAM_37 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_38 = 256'hFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00;
defparam sp_inst_7.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_3A = 256'hFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000F;
defparam sp_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_3C = 256'hF7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000FFFFFFFF;
defparam sp_inst_7.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7;
defparam sp_inst_7.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFF;
defparam sp_inst_7.INIT_RAM_3F = 256'hFFFFFFFFF7F7F7F00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F7F7F0000;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[29:0],sp_inst_8_dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b00;
defparam sp_inst_8.BIT_WIDTH = 2;
defparam sp_inst_8.BLK_SEL = 3'b010;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'h2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA;
defparam sp_inst_8.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFF;
defparam sp_inst_8.INIT_RAM_03 = 256'hC0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_04 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500;
defparam sp_inst_8.INIT_RAM_06 = 256'hFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_07 = 256'hAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2A;
defparam sp_inst_8.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFF;
defparam sp_inst_8.INIT_RAM_0A = 256'hFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF;
defparam sp_inst_8.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA155515550000;
defparam sp_inst_8.INIT_RAM_0D = 256'hFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_0E = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000;
defparam sp_inst_8.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_11 = 256'h3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_12 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF;
defparam sp_inst_8.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA15551555000000;
defparam sp_inst_8.INIT_RAM_14 = 256'hFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_15 = 256'h55155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA15;
defparam sp_inst_8.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_18 = 256'hFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3F;
defparam sp_inst_8.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000;
defparam sp_inst_8.INIT_RAM_1B = 256'hFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_1C = 256'h155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555;
defparam sp_inst_8.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_1F = 256'h2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF;
defparam sp_inst_8.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFF2AAA2AAA1555155500000000FF;
defparam sp_inst_8.INIT_RAM_22 = 256'hFFFFEFFF3FFF2AAA2AAA1555155500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_23 = 256'h5500000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAA2AAA15551555155515;
defparam sp_inst_8.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_28 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce_w)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_2_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(sp_inst_1_dout[1]),
  .I1(sp_inst_2_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(sp_inst_3_dout[2]),
  .I1(sp_inst_5_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(sp_inst_4_dout[3]),
  .I1(sp_inst_5_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(sp_inst_6_dout[4]),
  .I1(sp_inst_8_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(sp_inst_7_dout[5]),
  .I1(sp_inst_8_dout[5]),
  .S0(dff_q_0)
);
endmodule //sp_framebuffer
